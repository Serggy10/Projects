* C:\Users\sergi\OneDrive\Escritorio\Comedero\MSIM\prueba1.sch

* Schematics Version 8.0 - July 1997
* Sun Jul 17 18:54:53 2022



** Analysis setup **
.tran 20ns 4s
.OP 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib "u:\Userlib\DTE_DIGITAL.lib"
.lib "u:\UserLib\DTE_1.lib"
.lib "nom.lib"

.INC "prueba1.net"
.INC "prueba1.als"


.probe


.END
