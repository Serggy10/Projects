* C:\Users\sergi\OneDrive\Escritorio\Comedero\prueba_emergencia.sch

* Schematics Version 8.0 - July 1997
* Wed Jul 20 12:22:11 2022



** Analysis setup **
.tran 20ns 2s
.OP 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib "u:\Userlib\DTE_DIGITAL.lib"
.lib "u:\UserLib\DTE_1.lib"
.lib "nom.lib"

.INC "prueba_emergencia.net"
.INC "prueba_emergencia.als"


.probe


.END
